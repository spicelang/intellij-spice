f<int> main() {
    printf("test: %d", 1.0);
    char test = 'a';
}